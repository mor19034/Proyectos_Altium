* STD2NA60 model from ST Microelectronics

.SUBCKT std2na60 1 2 3
LG 2 4  7.5n
LS 12 3 7.5n
LD 6 1  4.5n
RG 4 5  2.05
RS 9 12 0.297383E-03
RD 7 6  2.83524
RJ 8 7  0.443553E-01
CGS 5 9  0.674320E-12
CGD 7 10 0.831998E-10
CK  11 7 0.131084E-10
DGD 11 7 DGD
DBS 12 6 DBS
DBD  9 7 DBD
MOS  13 5 9 9 MOS L=0.311893E-05 W=0.686489
E1  10 5 101 0 1
E2  11 5 102 0 1
E3  8 13 POLY(2) 6 8 6 12 0 0 0 0  0.338138E-01
G1  0 100 7 5 1u
D1  100 101  DID
D2  102 100  DID
R1  101 0  1MEG
R2  102 0  1MEG
.MODEL MOS NMOS
+ LEVEL = 3
+ TOX   = .11E-06
+ VTO   = 3.96762
+ PHI   = 1.68193
+ NSUB  = .52E+17
+ IS    = 0
+ JS    = 0
+ UO    = 420
+ THETA = .05
+ KP    = 0.146889E-04
.MODEL DGD D
+ CJO   =0.616243E-09
+ VJ    =0.454980
+ M     =0.744248
.MODEL DBD D
+ CJO   =0.347939E-09
+ VJ    =0.649211
+ M     =0.783001
.MODEL DBS D
+ IS    =0.1P
+ BV    = 661.902
+ N     = 1
+ TT    = .246679E-06
+ RS    =4.55M
.MODEL DID D
+ IS    =2P
+ RS    = 0
+ BV    = 671.902
.ENDS std2na60

