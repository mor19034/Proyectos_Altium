**********
*==========================================================
* UC3842B
* ON Semiconductor
* PWM Controller
*
* This model was developed for ON Semiconductor by:
* AEI Systems, LLC
* 5777 W. Century Blvd. Suite 876
* Los Angeles, California 90045
* Copyright 2002, all rights reserved.
*
* This model is subject to change without notice.
* Users may not directly or indirectly re-sell or
* re-distribute this model. This model may not
* be used, modified, or altered
* without the consent of ON Semiconductor.
*
* For more information regarding modeling services,
* model libraries and simulation products, please
* call AEi Systems at (310) 863-8034, or contact
* AEi by email: info@aeng.com. http://www.AENG.com
*
* Revision: 1.0
*==========================================================
* CLS translated PSpice syntax to XSpice
*SRC=UC3842B;UC3842B;ON Semiconductor;PWM Controllers;96% DC, 16V/10V
*SYM=UC3845
.SUBCKT UC3842B  3    14   15   1     18    4   20   2
*              E/A  FDBK  IS  RT/CT  GND  OUT  VC  VREF
*
.SUBCKT 1845AMP  4     1    9   20
*                VREF  INV  OUT V-
.MODEL QPMOD PNP
.MODEL DCLAMP D (RS=10 BV=5 IBV=.01)
.MODEL DMOD D
R1 10 4 100K
R2 10 20 100K
R3 6 20 316MEG
C1 6 20 15.9P
E1 5 20 6 20 1
R4 1 20 8MEG
I2 4 9 .8M
D12 9 4 DMOD
R6 20 3 300
D11 9 12 DMOD
Q1 20 13 12 QPMOD
I3 13 20 68U
D14 3 13 DMOD
D15 20 6 DCLAMP
L1 2 3 10U
C2 3 20 200P
R9 5 2 5
C5 2 20 .02U
G1 20 6 10 1 100U
.ENDS
*
.SUBCKT 1845OUT  4  7  3  12
*                +V -V IN OUT
.MODEL QMOD NPN RC=1.5 RE=.5 RB=100 IKF=0.5 CJC=0.4P
.MODEL QMOD2 NPN TF=400P TR=400P
.MODEL QIN NPN BF=100 BR=2 IS=1E-16 VAF=50 
+ CJE=1.5P CJC=.15P TR=1N TF=4N
.MODEL DMOD D RS=1 IS=0.4U
I3 4 8 100U
D3 8 4 DMOD
D4 12 8 DMOD
Q3 8 1 9 QIN
Q4 12 9 7 QMOD
Q5 4 8 6 QMOD
I4 7 1 .9M
R1 3 2 10K
Q8 1 2 7 QIN
Q2 4 6 12 QMOD2
.ENDS
*
.SUBCKT FFLOP     1    2  11 12  5     6
*                 CLK  D  R  S   QBAR  Q
.SUBCKT NAND3 1 2 3 4 params: IC=0
B1 5 0 V=~(V(1)&V(2)&V(3))
R1 5 4 400
C1 4 0 20P IC={IC}
.ENDS
.SUBCKT INV 1 2 params: IC=0
B1 3 0 V=~(V(1))
R1 3 2 100
C1 2 0 10P IC={IC}
.ENDS
X1 7 4 2 8 NAND3 params: IC=0
X2 8 3 10 9 NAND3 params: IC=0
X3 1 8 10 7 NAND3 params: IC=3.5
X4 4 9 1 10 NAND3 params: IC=0
X5 4 7 6 5 NAND3 params: IC=3.5
X6 5 10 3 6 NAND3 params: IC=0
X7 11 4 INV params: IC=3.5
X8 12 3 INV params: IC=3.5
.ENDS
*
****OSCILLATOR*****
S1 8 18 1 18 SOSC
.MODEL SOSC SW(RON=.01 ROFF=1MEG VT=2.05 VH=.8)
BDISCH 1 18 I=8.3m * u(2.5-V(8,18)) * u(V(13,18)-2.5)
RPULL 8 2 100K
****UVLO***********
S4 20 19 20 18 SUVLO
.MODEL SUVLO SW(RON=.01 ROFF=1MEG VT=13 VH=3)
RUVLO 19 18 1MEG
RSTDBY 20 18 32K
ROP 10 18 500
****REFERENCE*******
BREF 13 18 V=5*u(V(19,18)-6)
RREG 10 2 .33
CREF 2 18 1n
V3 13 10 0V
B6 19 18 I=I(V3)
****CURRENT COMPARATOR*******
B3 21 18 V=5*u(V(15,18) - V(16,18))
R7 15 18 1MEG
RDELAY 21 22 1K
CDELAY 22 18 150P
****ERROR AMPLIFIER**********
XAMP 2 14 3 18 1845AMP
****OFFSET LIMITER***********
R4 12 11 2MEG
R6 11 18 1MEG
B2 16 18 V=1 - uramp(1-V(11,18))
V4 3 9 1
D1 9 12 D2
.MODEL D2 D 
****OUTPUT DRIVER************
XDRIVE 19 18 5 4 1845OUT
****S-R LATCH****************
XLATCH 8 2 22 18 6 7 FFLOP params: 
****OUTPUT AND GATE**********
B8 5 18 V=10 * u(V(2,18)-2.5) * u(V(7,18)-2.5) *u(V(8,18)-2.5)
.ENDS
