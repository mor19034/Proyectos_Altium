*Simplified Transformer Subcircuit Parameters
*L1     = primary inductance
*RATIO1 = turns ratio (= secondary1/primary)
*RATIO2 = turns ratio (= secondary2/primary)
*
*Connections:
*                    Pri+
*                    | Pri-
*                    | | Sec1+
*                    | | | Sec1-
*                    | | | | Sec2+
*                    | | | | | Sec2-
*                    | | | | | |
.SUBCKT SIMPL3WTRANS 1 2 3 4 5 6 PARAMS: L1=1m RATIO1=1 RATIO2=1
Lx 1 2 {L1}
Xx 1 2 3 4 5 6 IDEAL3W PARAMS: RATIO1={RATIO1} RATIO2={RATIO2}
.SUBCKT IDEAL3W 1 2 3 4 5 6 PARAMS: RATIO1=1 RATIO2=1
BP  1 2 I=( -I(BS1)*{RATIO1} - I(BS2)*{RATIO2} )
BS1 3 4 V=( V(1,2)*{RATIO1} )
BS2 5 6 V=( V(1,2)*{RATIO2} )
.ENDS IDEAL3W
.ENDS SIMPL3WTRANS
