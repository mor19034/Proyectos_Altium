* General-purpose optocoupler model derived from Transim circuit templates

.SUBCKT GEN_OPTO A K C E
C1   6 K 4u
D1   A 5 IDEAL
.MODEL IDEAL D(IS=1p)
F1   K 6 VF1 2
VF1  5 K 0
G1   C E 6 K 1
R1   6 K 1
X$R2 E C SIMPLIS_VPWLR_R2 PARAMS: IC=1
.SUBCKT SIMPLIS_VPWLR_R2 1 2 PARAMS: IC=1 NSEG=3 X0=-100 Y0=-1e-6 X1=0.00 Y1=0 X2=.001 Y2=1e-3 X3=0.01 Y3=1
.PARAM C = {(X1*Y0 - X0*Y1) / (X1 - X0)}
.PARAM A0 = {(Y1 - Y0) / (X1 - X0)}
.PARAM A1 = {(Y2 - Y1) / (X2 - X1) - A0}
.PARAM A2 = {(Y3 - Y2) / (X3 - X2) - A0 - A1}
Bx 1 2 I = C + A0*v(1,2) + A1*uramp(v(1,2)-X1) + A2*uramp(v(1,2)-X2)
.ENDS SIMPLIS_VPWLR_R2
.ENDS GEN_OPTO
